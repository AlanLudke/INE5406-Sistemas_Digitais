#�d�(��oh	�|�rַ���_u��}�J�5�e�3Z�%y��0v�;@�dC��NCx�F$Ș�h��#�T�,O�(�C��4o"�wQ(�W���2u��M���E����ӱR{���2
%/�kL� ��`j��Gc�Y̩_����@�^�9X�my��`X�5�&0�0$_�*5��b��)"<oS�R�|ϭ[4R �4���g8�۟�c�I*dT!}0��g��K�{ �{��?H-��,��T�%���U�8�O�;�w��Gu)���ؑ�S{m��^ v�=F�����Q��bli����0S�a� y�2C�0P�@; �e#d�#���#|1>
odF��^�3�/�YM�2��g���GђW� �l�<)�*���}y�>��#_��{�o|G?	���x
��@�$��g4�0����*�}tr	x�T��Ȇn�|�-�G�P$��'��^��Zuv�sl���K?�d`�r����{�y����eS��ٸ���oA���'[#��Գ����$M�ӳ���p0�ަ�:�Y�-���$�6��M�b��Y�v3�U��9C"A��6��k�m�8��8 3^��,��H�%$p�)͢૰G�W�O�����o��"/�%3�x#�,���I��a�lV�r��m�t)aj�$\��xM��K��=���L�D�����"��٦�ǋ�ظ��%O�3d�lk-��]8��R��%KԖ�#ڽ��E�V_h���g�bz2���H�w�GD�m�o3v��Qj�����	��������;��J�R��-���i�d�z��\��:�ԃ� ܌�B4D@�HM�[��Skz�gs��O��W(ϯ����=^p���N@�O��j�-��f"C�wR��1`��ۻ�_/�$�$Xi9dM��L��NZ3_���u�v��뮽w��s�bXe�T��R:�g��a�!�5 LJ������"�f�5