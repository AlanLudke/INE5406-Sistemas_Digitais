����vU}�������=}[�3;w�ҵ��RM�Vw�?ͭ+P��ާ��M�ӱ���	9�����֢[��+1��a���]�!� A�d�bwo�G�f���&ؚ���$W����v|N�.��1*&b0jt��ό�Z��Q�X�
�r)�1�v��m���l&wlလ�
�m�y��.֬���1e�,/q�R3H-N��\Z}�ى8�#�۩Xs>�_ ��Ҥ�X��Ud�L�F���C|S&��>�^�W|CR��1���DWQ�耣�ū\���Nu�X��M������ݒݷ�t=ׂ�o0�<#������iA"K�V*�6h�]�!l�ǷNge�N�z>������r�H�j�r�~{*㭡�����ݱ��k�;zof�,��Fk�8��;<<����E�
t���	$���$ϗjZ�.%mNhM��R��������981(T���׺�Q-���#	�Xܼѥ{*5l�;�BŜ!�>6_���� �/0��YPO���w�d�N�=�~�K���l��Mtw����XX��dC��.��9��6��w��z�8J):�rIA��X$�G��0�
3��#��1rA#';"�o�?���%&M����$�U��I��e��OKYc���krw_}E/�\7��k�W���˴���i�`���3ְO%�/UjU��6n�1����LT��U����'i˵���<�