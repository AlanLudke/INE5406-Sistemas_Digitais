� r�U��f'�^�
��,��h��Kp����d���z��VpܬD�����<�N��	I���f���f��e�@u�\��z��4�>��x��|�`\�@��7�I�j�g8�$����\��8�}�xZ��+@	S7��(���4؏_��^�J����?�-�y�]���j���n��n������4�'��Z��@��B��;.�ċ�0+����H,*�T4��a��,{�w�ɨ�^��텺�4�̲�5�*��_�ǃɔ/��T�����01c�y�{տG�<t#i�^�B�lA*78�gq=��|d:�/�	g'��N^8�`��0�A�3�ł6lI��5���t�M؃�H wY[|��]�������k7�d���M��W[�;J�T�>FA;Q@0nC�I�AJ����!�i)������D��=��,����7����/�S�ߺb�)�޻|Vaa���zn�~k�*�y�yKj}�PRBL���K�0�����:;�·+e (hW<��iY��{y��;�Ԕ�)p���G[?"0iTJܯ�(�ugA��q��ٜ�	os�F]\�,zP����8�#f��-C��Y`��s)��K<�)�0�}9�K��]s�B"-b,|'�d��w� Wa��x;��߸�o���V"iRj��W���*���5�T��KrY�Y�����Jkv0��=�!�����D{����L���G\�%KlE5}d/.�s��ߖ��Cٯ�����%�"����zj�Ca��rn�A�C�s¢:̜B�s҆G�	��|�FP��9@I�?���o.ݯ����RGBi6ӸTDG3�&�J:��P�����04 �B�YpXգ
��n�LULob�L���/��P��xu�پ�g$Xq��^L0�F�ψ�j����� R��77�^h�I]��Ys=х���'�o�o�����!��wτ�1;xͤ�Zm���bj����m�ݔ�h��o@<�^k)���8M*E�<�zk��7�koh����s�}�lw6���\kY�I[p+�"�G�é�����(�)����=��vk{��(���4�{�7H��x5� ����g��=6|5�}